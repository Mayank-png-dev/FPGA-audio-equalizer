//fft_1024.v
module fft_1024
    input clk,
    input rst,
    input signed [15:0] data_in,
    input data_valid,
    output signed [15:0] data_out_real,
    output signed [15:0] data_out_imag,
    output out_valid
);
    // T0Do: Implement radix-2 fft
endmodule